library ieee;
use ieee.std_logic_1164.all;
use work.system_components.all;

entity phase1 is
	port (
		R : in std_logic -- to be replaced later on with proper ports
	);
end entity;

architecture arch_phase1 of phase1 is

begin

end architecture;