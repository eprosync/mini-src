// welcome to my personal hell.
// this is for the final project, phase4.
module computer()

endmodule