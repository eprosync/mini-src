module op_shla_32(input [31:0] Ain, Bin, output [31:0] Zout);
    assign Zout = $signed(Ain) << Bin;
endmodule