-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Mon Feb 13 16:35:43 2023"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY alu IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		CS :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		C :  OUT  STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END alu;

ARCHITECTURE bdf_type OF alu IS 

COMPONENT alu_32_to_64
	PORT(en : IN STD_LOGIC;
		 C_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C_in_64 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 C_out : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_divide0
	PORT(denom : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 numer : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 quotient : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 remain : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_add_32
	PORT(Cin : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Cout : OUT STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu_guard_switch
	PORT(en : IN STD_LOGIC;
		 A_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 A_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_and_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu_op_combiner
	PORT(op_add_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_and_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_div_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_mul_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_negate_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_not_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_or_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_rol_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_ror_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_shl_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_shr_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 op_sub_in : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 C_out : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu_op_decider
	PORT(CS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 op_add : OUT STD_LOGIC;
		 op_sub : OUT STD_LOGIC;
		 op_mul : OUT STD_LOGIC;
		 op_div : OUT STD_LOGIC;
		 op_and : OUT STD_LOGIC;
		 op_or : OUT STD_LOGIC;
		 op_shr : OUT STD_LOGIC;
		 op_shl : OUT STD_LOGIC;
		 op_ror : OUT STD_LOGIC;
		 op_rol : OUT STD_LOGIC;
		 op_not : OUT STD_LOGIC;
		 op_negate : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT op_mul_32
	PORT(M : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Q : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 P : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_not_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_or_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_rol_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_ror_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_shl_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT op_shr_32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 C : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(0 TO 63);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC_VECTOR(31 DOWNTO 0);


BEGIN 
SYNTHESIZED_WIRE_2 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_5 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_8 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_11 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_14 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_18 <= "00000000000000000000000000000000";
SYNTHESIZED_WIRE_22 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_25 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_28 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_31 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_34 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_37 <= "0000000000000000000000000000000000000000000000000000000000000000";
SYNTHESIZED_WIRE_38 <= '0';
SYNTHESIZED_WIRE_61 <= '1';
SYNTHESIZED_WIRE_63 <= "00000000000000000000000000000000";
SYNTHESIZED_WIRE_83 <= '1';
SYNTHESIZED_WIRE_85 <= "00000000000000000000000000000000";
SYNTHESIZED_WIRE_86 <= '0';



b2v_inst : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_91,
		 C_in => SYNTHESIZED_WIRE_1,
		 C_in_64 => SYNTHESIZED_WIRE_2,
		 C_out => SYNTHESIZED_WIRE_45);


b2v_inst1 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_92,
		 C_in => SYNTHESIZED_WIRE_4,
		 C_in_64 => SYNTHESIZED_WIRE_5,
		 C_out => SYNTHESIZED_WIRE_56);


b2v_inst10 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_93,
		 C_in => SYNTHESIZED_WIRE_7,
		 C_in_64 => SYNTHESIZED_WIRE_8,
		 C_out => SYNTHESIZED_WIRE_52);


b2v_inst11 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_94,
		 C_in => SYNTHESIZED_WIRE_10,
		 C_in_64 => SYNTHESIZED_WIRE_11,
		 C_out => SYNTHESIZED_WIRE_50);


b2v_inst12 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_95,
		 C_in => SYNTHESIZED_WIRE_13,
		 C_in_64 => SYNTHESIZED_WIRE_14,
		 C_out => SYNTHESIZED_WIRE_49);


b2v_inst14 : lpm_divide0
PORT MAP(denom => SYNTHESIZED_WIRE_15,
		 numer => SYNTHESIZED_WIRE_16,
		 quotient => SYNTHESIZED_WIRE_21);


b2v_inst2 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_96,
		 C_in => SYNTHESIZED_WIRE_18,
		 C_in_64 => SYNTHESIZED_WIRE_19,
		 C_out => SYNTHESIZED_WIRE_48);










b2v_inst4 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_97,
		 C_in => SYNTHESIZED_WIRE_21,
		 C_in_64 => SYNTHESIZED_WIRE_22,
		 C_out => SYNTHESIZED_WIRE_47);












b2v_inst5 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_98,
		 C_in => SYNTHESIZED_WIRE_24,
		 C_in_64 => SYNTHESIZED_WIRE_25,
		 C_out => SYNTHESIZED_WIRE_46);


b2v_inst6 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_99,
		 C_in => SYNTHESIZED_WIRE_27,
		 C_in_64 => SYNTHESIZED_WIRE_28,
		 C_out => SYNTHESIZED_WIRE_51);


b2v_inst7 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_100,
		 C_in => SYNTHESIZED_WIRE_30,
		 C_in_64 => SYNTHESIZED_WIRE_31,
		 C_out => SYNTHESIZED_WIRE_55);


b2v_inst8 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_101,
		 C_in => SYNTHESIZED_WIRE_33,
		 C_in_64 => SYNTHESIZED_WIRE_34,
		 C_out => SYNTHESIZED_WIRE_54);


b2v_inst9 : alu_32_to_64
PORT MAP(en => SYNTHESIZED_WIRE_102,
		 C_in => SYNTHESIZED_WIRE_36,
		 C_in_64 => SYNTHESIZED_WIRE_37,
		 C_out => SYNTHESIZED_WIRE_53);


b2v_op_add : op_add_32
PORT MAP(Cin => SYNTHESIZED_WIRE_38,
		 A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_40,
		 S => SYNTHESIZED_WIRE_1);


b2v_op_add_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_91,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_39,
		 B_out => SYNTHESIZED_WIRE_40);


b2v_op_and : op_and_32
PORT MAP(A => SYNTHESIZED_WIRE_42,
		 B => SYNTHESIZED_WIRE_43,
		 C => SYNTHESIZED_WIRE_24);


b2v_op_and_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_98,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_42,
		 B_out => SYNTHESIZED_WIRE_43);


b2v_op_combiner : alu_op_combiner
PORT MAP(op_add_in => SYNTHESIZED_WIRE_45,
		 op_and_in => SYNTHESIZED_WIRE_46,
		 op_div_in => SYNTHESIZED_WIRE_47,
		 op_mul_in => SYNTHESIZED_WIRE_48,
		 op_negate_in => SYNTHESIZED_WIRE_49,
		 op_not_in => SYNTHESIZED_WIRE_50,
		 op_or_in => SYNTHESIZED_WIRE_51,
		 op_rol_in => SYNTHESIZED_WIRE_52,
		 op_ror_in => SYNTHESIZED_WIRE_53,
		 op_shl_in => SYNTHESIZED_WIRE_54,
		 op_shr_in => SYNTHESIZED_WIRE_55,
		 op_sub_in => SYNTHESIZED_WIRE_56,
		 C_out => C);


b2v_op_decider : alu_op_decider
PORT MAP(CS => CS,
		 op_add => SYNTHESIZED_WIRE_91,
		 op_sub => SYNTHESIZED_WIRE_92,
		 op_mul => SYNTHESIZED_WIRE_96,
		 op_div => SYNTHESIZED_WIRE_97,
		 op_and => SYNTHESIZED_WIRE_98,
		 op_or => SYNTHESIZED_WIRE_99,
		 op_shr => SYNTHESIZED_WIRE_100,
		 op_shl => SYNTHESIZED_WIRE_101,
		 op_ror => SYNTHESIZED_WIRE_102,
		 op_rol => SYNTHESIZED_WIRE_93,
		 op_not => SYNTHESIZED_WIRE_94,
		 op_negate => SYNTHESIZED_WIRE_95);


b2v_op_divide_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_97,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_16,
		 B_out => SYNTHESIZED_WIRE_15);


b2v_op_mul : op_mul_32
PORT MAP(M => SYNTHESIZED_WIRE_58,
		 Q => SYNTHESIZED_WIRE_59,
		 P => SYNTHESIZED_WIRE_19);


b2v_op_mul_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_96,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_58,
		 B_out => SYNTHESIZED_WIRE_59);


b2v_op_negate_2s_comp : op_add_32
PORT MAP(Cin => SYNTHESIZED_WIRE_61,
		 A => SYNTHESIZED_WIRE_62,
		 B => SYNTHESIZED_WIRE_63,
		 S => SYNTHESIZED_WIRE_13);


b2v_op_negate_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_95,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_65);


b2v_op_negate_not : op_not_32
PORT MAP(A => SYNTHESIZED_WIRE_65,
		 C => SYNTHESIZED_WIRE_62);


b2v_op_not : op_not_32
PORT MAP(A => SYNTHESIZED_WIRE_66,
		 C => SYNTHESIZED_WIRE_10);


b2v_op_not_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_94,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_66);


b2v_op_or : op_or_32
PORT MAP(A => SYNTHESIZED_WIRE_68,
		 B => SYNTHESIZED_WIRE_69,
		 C => SYNTHESIZED_WIRE_27);


b2v_op_or_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_99,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_68,
		 B_out => SYNTHESIZED_WIRE_69);


b2v_op_rol : op_rol_32
PORT MAP(A => SYNTHESIZED_WIRE_71,
		 B => SYNTHESIZED_WIRE_72,
		 C => SYNTHESIZED_WIRE_7);


b2v_op_rol_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_93,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_71,
		 B_out => SYNTHESIZED_WIRE_72);


b2v_op_ror : op_ror_32
PORT MAP(A => SYNTHESIZED_WIRE_74,
		 B => SYNTHESIZED_WIRE_75,
		 C => SYNTHESIZED_WIRE_36);


b2v_op_ror_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_102,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_74,
		 B_out => SYNTHESIZED_WIRE_75);


b2v_op_shl : op_shl_32
PORT MAP(A => SYNTHESIZED_WIRE_77,
		 B => SYNTHESIZED_WIRE_78,
		 C => SYNTHESIZED_WIRE_33);


b2v_op_shl_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_101,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_77,
		 B_out => SYNTHESIZED_WIRE_78);


b2v_op_shr : op_shr_32
PORT MAP(A => SYNTHESIZED_WIRE_80,
		 B => SYNTHESIZED_WIRE_81,
		 C => SYNTHESIZED_WIRE_30);


b2v_op_shr_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_100,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_80,
		 B_out => SYNTHESIZED_WIRE_81);


b2v_op_sub_2s_comp : op_add_32
PORT MAP(Cin => SYNTHESIZED_WIRE_83,
		 A => SYNTHESIZED_WIRE_84,
		 B => SYNTHESIZED_WIRE_85,
		 S => SYNTHESIZED_WIRE_88);


b2v_op_sub_adder : op_add_32
PORT MAP(Cin => SYNTHESIZED_WIRE_86,
		 A => SYNTHESIZED_WIRE_87,
		 B => SYNTHESIZED_WIRE_88,
		 S => SYNTHESIZED_WIRE_4);


b2v_op_sub_guard : alu_guard_switch
PORT MAP(en => SYNTHESIZED_WIRE_92,
		 A_in => A,
		 B_in => B,
		 A_out => SYNTHESIZED_WIRE_87,
		 B_out => SYNTHESIZED_WIRE_90);


b2v_op_sub_invert : op_not_32
PORT MAP(A => SYNTHESIZED_WIRE_90,
		 C => SYNTHESIZED_WIRE_84);


END bdf_type;