library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.system_components.all;

entity ALU_tb is
	
end;

architecture ALU_tb_behavioral of ALU_tb is

begin

end architecture;